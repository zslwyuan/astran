.subckt AND2X1INV Q B VCC GND A
M0 a_2_6# A VCC VCC PMOS L=65n W=500n
M1 VCC B a_2_6# VCC PMOS L=65n W=500n
M2 Y a_2_6# VCC VCC PMOS L=65n W=500n
M3 a_9_6# A a_2_6# GND NMOS L=65n W=500n
M4 GND B a_9_6# GND NMOS L=65n W=500n
M5 Y a_2_6# GND GND NMOS L=65n W=500n
MN Q Y GND GND nmos L=65n W=240n
MP Q Y VCC VCC pmos L=65n W=520n
.ends

